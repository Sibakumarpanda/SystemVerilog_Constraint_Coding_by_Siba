//21.WAC to generate Even numbers in odd positions and a value of 50 in all even positions with in range 1-100

class my_packet;
  rand int a [];
  //rand bit a [];  
  //constraint c1 {a inside {[1:100]};}  
  constraint c1 {a.size == 100;}
  constraint c2 { foreach (a[i])
                     if (i%2 !=0)
                       a[i] == i+1; // At Odd Positions
                     else
                       a[i] == 50 ; //At all Even Positions , value should be 50                                            
                }  
endclass 

module tb_top;  
  initial begin   
    my_packet pkt;
    pkt=new();    
    for (int i=0; i<10;i++) begin
      pkt.randomize();
      $display("The Generated Pattern in %0d iteration : a=%p",i,pkt.a); 
    end 
  end  
endmodule  
//output
The Generated Pattern in 0 iteration : a='{50, 2, 50, 4, 50, 6, 50, 8, 50, 10, 50, 12, 50, 14, 50, 16, 50, 18, 50, 20, 50, 22, 50, 24, 50, 26, 50, 28, 50, 30, 50, 32, 50, 34, 50, 36, 50, 38, 50, 40, 50, 42, 50, 44, 50, 46, 50, 48, 50, 50, 50, 52, 50, 54, 50, 56, 50, 58, 50, 60, 50, 62, 50, 64, 50, 66, 50, 68, 50, 70, 50, 72, 50, 74, 50, 76, 50, 78, 50, 80, 50, 82, 50, 84, 50, 86, 50, 88, 50, 90, 50, 92, 50, 94, 50, 96, 50, 98, 50, 100} 
The Generated Pattern in 1 iteration : a='{50, 2, 50, 4, 50, 6, 50, 8, 50, 10, 50, 12, 50, 14, 50, 16, 50, 18, 50, 20, 50, 22, 50, 24, 50, 26, 50, 28, 50, 30, 50, 32, 50, 34, 50, 36, 50, 38, 50, 40, 50, 42, 50, 44, 50, 46, 50, 48, 50, 50, 50, 52, 50, 54, 50, 56, 50, 58, 50, 60, 50, 62, 50, 64, 50, 66, 50, 68, 50, 70, 50, 72, 50, 74, 50, 76, 50, 78, 50, 80, 50, 82, 50, 84, 50, 86, 50, 88, 50, 90, 50, 92, 50, 94, 50, 96, 50, 98, 50, 100} 
The Generated Pattern in 2 iteration : a='{50, 2, 50, 4, 50, 6, 50, 8, 50, 10, 50, 12, 50, 14, 50, 16, 50, 18, 50, 20, 50, 22, 50, 24, 50, 26, 50, 28, 50, 30, 50, 32, 50, 34, 50, 36, 50, 38, 50, 40, 50, 42, 50, 44, 50, 46, 50, 48, 50, 50, 50, 52, 50, 54, 50, 56, 50, 58, 50, 60, 50, 62, 50, 64, 50, 66, 50, 68, 50, 70, 50, 72, 50, 74, 50, 76, 50, 78, 50, 80, 50, 82, 50, 84, 50, 86, 50, 88, 50, 90, 50, 92, 50, 94, 50, 96, 50, 98, 50, 100} 
The Generated Pattern in 3 iteration : a='{50, 2, 50, 4, 50, 6, 50, 8, 50, 10, 50, 12, 50, 14, 50, 16, 50, 18, 50, 20, 50, 22, 50, 24, 50, 26, 50, 28, 50, 30, 50, 32, 50, 34, 50, 36, 50, 38, 50, 40, 50, 42, 50, 44, 50, 46, 50, 48, 50, 50, 50, 52, 50, 54, 50, 56, 50, 58, 50, 60, 50, 62, 50, 64, 50, 66, 50, 68, 50, 70, 50, 72, 50, 74, 50, 76, 50, 78, 50, 80, 50, 82, 50, 84, 50, 86, 50, 88, 50, 90, 50, 92, 50, 94, 50, 96, 50, 98, 50, 100} 
The Generated Pattern in 4 iteration : a='{50, 2, 50, 4, 50, 6, 50, 8, 50, 10, 50, 12, 50, 14, 50, 16, 50, 18, 50, 20, 50, 22, 50, 24, 50, 26, 50, 28, 50, 30, 50, 32, 50, 34, 50, 36, 50, 38, 50, 40, 50, 42, 50, 44, 50, 46, 50, 48, 50, 50, 50, 52, 50, 54, 50, 56, 50, 58, 50, 60, 50, 62, 50, 64, 50, 66, 50, 68, 50, 70, 50, 72, 50, 74, 50, 76, 50, 78, 50, 80, 50, 82, 50, 84, 50, 86, 50, 88, 50, 90, 50, 92, 50, 94, 50, 96, 50, 98, 50, 100} 
The Generated Pattern in 5 iteration : a='{50, 2, 50, 4, 50, 6, 50, 8, 50, 10, 50, 12, 50, 14, 50, 16, 50, 18, 50, 20, 50, 22, 50, 24, 50, 26, 50, 28, 50, 30, 50, 32, 50, 34, 50, 36, 50, 38, 50, 40, 50, 42, 50, 44, 50, 46, 50, 48, 50, 50, 50, 52, 50, 54, 50, 56, 50, 58, 50, 60, 50, 62, 50, 64, 50, 66, 50, 68, 50, 70, 50, 72, 50, 74, 50, 76, 50, 78, 50, 80, 50, 82, 50, 84, 50, 86, 50, 88, 50, 90, 50, 92, 50, 94, 50, 96, 50, 98, 50, 100} 
The Generated Pattern in 6 iteration : a='{50, 2, 50, 4, 50, 6, 50, 8, 50, 10, 50, 12, 50, 14, 50, 16, 50, 18, 50, 20, 50, 22, 50, 24, 50, 26, 50, 28, 50, 30, 50, 32, 50, 34, 50, 36, 50, 38, 50, 40, 50, 42, 50, 44, 50, 46, 50, 48, 50, 50, 50, 52, 50, 54, 50, 56, 50, 58, 50, 60, 50, 62, 50, 64, 50, 66, 50, 68, 50, 70, 50, 72, 50, 74, 50, 76, 50, 78, 50, 80, 50, 82, 50, 84, 50, 86, 50, 88, 50, 90, 50, 92, 50, 94, 50, 96, 50, 98, 50, 100} 
The Generated Pattern in 7 iteration : a='{50, 2, 50, 4, 50, 6, 50, 8, 50, 10, 50, 12, 50, 14, 50, 16, 50, 18, 50, 20, 50, 22, 50, 24, 50, 26, 50, 28, 50, 30, 50, 32, 50, 34, 50, 36, 50, 38, 50, 40, 50, 42, 50, 44, 50, 46, 50, 48, 50, 50, 50, 52, 50, 54, 50, 56, 50, 58, 50, 60, 50, 62, 50, 64, 50, 66, 50, 68, 50, 70, 50, 72, 50, 74, 50, 76, 50, 78, 50, 80, 50, 82, 50, 84, 50, 86, 50, 88, 50, 90, 50, 92, 50, 94, 50, 96, 50, 98, 50, 100} 
The Generated Pattern in 8 iteration : a='{50, 2, 50, 4, 50, 6, 50, 8, 50, 10, 50, 12, 50, 14, 50, 16, 50, 18, 50, 20, 50, 22, 50, 24, 50, 26, 50, 28, 50, 30, 50, 32, 50, 34, 50, 36, 50, 38, 50, 40, 50, 42, 50, 44, 50, 46, 50, 48, 50, 50, 50, 52, 50, 54, 50, 56, 50, 58, 50, 60, 50, 62, 50, 64, 50, 66, 50, 68, 50, 70, 50, 72, 50, 74, 50, 76, 50, 78, 50, 80, 50, 82, 50, 84, 50, 86, 50, 88, 50, 90, 50, 92, 50, 94, 50, 96, 50, 98, 50, 100} 
The Generated Pattern in 9 iteration : a='{50, 2, 50, 4, 50, 6, 50, 8, 50, 10, 50, 12, 50, 14, 50, 16, 50, 18, 50, 20, 50, 22, 50, 24, 50, 26, 50, 28, 50, 30, 50, 32, 50, 34, 50, 36, 50, 38, 50, 40, 50, 42, 50, 44, 50, 46, 50, 48, 50, 50, 50, 52, 50, 54, 50, 56, 50, 58, 50, 60, 50, 62, 50, 64, 50, 66, 50, 68, 50, 70, 50, 72, 50, 74, 50, 76, 50, 78, 50, 80, 50, 82, 50, 84, 50, 86, 50, 88, 50, 90, 50, 92, 50, 94, 50, 96, 50, 98, 50, 100} 
           V C S   S i m u l a t i o n   R e p o r t 
